module mini_counter(
input clk,
rst,
output reg [31:0] cnt
);



endmodule